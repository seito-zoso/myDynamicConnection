import( <cygwin_kernel.cdl> );

signature sDynamic {
    void say_str( void );
};
signature sGetDescriptor {
    void getDescriptor( [out] Descriptor(sDynamic) *pDesc, [in] int ith );
};

celltype tTaskMain {
    entry sTaskBody eBody;
    [dynamic, optional]
        call sDynamic cDynamic;
    [ref_desc, optional]
        call sDynamic cRefDesc[];
    call sGetDescriptor cGetDescriptor;
};

celltype tRefDesc {
    entry sGetDescriptor eGetDescriptor;
    [ref_desc, optional]
        call sDynamic cRefDesc[];
};

celltype tDynamic {
    entry sDynamic eDynamic;
    attr {
        char *str;
    };
};

/* 組み上げ */
cell tTask Task {
    taskAttribute = C_EXP("TA_ACT");
    priority      = 11;
    stackSize     = 4096;
    cBody         = rTEMP::TaskMain.eBody;
};

[in_through()] // リージョン内への結合の許可
region rTEMP {
    cell tTaskMain TaskMain {
        cGetDescriptor = RefDesc.eGetDescriptor;
        cRefDesc[] = DynamicA.eDynamic;
        cRefDesc[] = DynamicB.eDynamic;
    };
    cell tRefDesc RefDesc {
        cRefDesc[] = DynamicA.eDynamic;
        cRefDesc[] = DynamicB.eDynamic;
    };
    cell tDynamic DynamicA {
        str = "Hello A";
    };
    cell tDynamic DynamicB {
        str = "Hello B";
    };
};
