import( <cygwin_kernel.cdl> );
import( <TECSInfo.cdl> );
import( <TECSInfoAccessor.cdl> );
import( "HelloWorld.cdl" );

/*
 * TECSInfo 使用サンプル
 */

signature sDynamic {
    initialize();
    do_something();
    finalize();
};

signature sGetDescriptor {
    ER getDescriptor( [out] Descriptor(sDynamic) *pDesc );
};
signature sSetDescriptor {
    ER setDescriptor( [in] Descriptor(sDynamic) desc );
};

celltype tTaskMain {
    entry sTaskBody eBody;
    [dynamic]
        call sDynamic cDynamic;
    [ref_desc]
        call sDynamic cRefDesc;
    call sGetDescriptor cGetDescriptor;
    entry sSetDescriptor eSetDescriptor;
};

celltype tDynamic {
    entry sDynamic eDynamic;
};

cell tTask Task {
    taskAttribute = C_EXP("TA_ACT");
    priority      = 11;
    stackSize     = 4096;
    cBody         = rTEMP::TaskMain.eBody;
};

[in_through()] // リージョン内への結合の許可
region rTEMP{
    cell tTaskMain TaskMain {
        cTECSInfo  = TECSInfo.eTECSInfo;
    };

};
